-- Datapath
