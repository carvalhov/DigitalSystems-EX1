-- Controlador
