library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity comparador8b is
port (
      -- Port inputs
      clock     : in std_logic; 
      EntA,EntB : in std_logic_vector(7 downto 0); 
      -- Port Output
      Output    : out std_logic -- Output = 1 when A >= B else 0
 );
end comparador8b;
  
architecture Behavioral of comparador8b is

  
end Behavioral;
